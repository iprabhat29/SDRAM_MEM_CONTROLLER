module monitor(ddr_interface.MONITOR inf);
/*  initial begin
    $dumpfile("dump.vcd");
    $dumpvars(1);
  end*/
endmodule